module  RAM(	input CLOCK,
					input [16:0] CoverPixel,
					input [12:0] PlayPausePixel,
					input [13:0] TitlePixel,
					input [11:0] SpeedPixel,
					input SecondSong,RW,
		
		output logic [3:0] CoverArtColor,
		output logic [23:0] TitleColor, PlayPauseColor, SpeedColor
);

// mem has width of 3 bits and a total of 400 addresses
logic [3:0] GrenadeArtmem [0:89999];
logic [3:0] JustArtmem [0:89999];
logic [23:0] Speedmem [0:2499];
logic [23:0] Pausemem [0:5183];
logic [23:0] Playmem [0:5183];
logic [23:0] Titlemem [0:14999];
logic [23:0] Title2mem [0:14999];

initial
begin
	 $readmemh("CoverArt/GrenadeP.txt", GrenadeArtmem);
	 $readmemh("CoverArt/JustTheWayYouAre.txt", JustArtmem);
	 $readmemh("CoverArt/icon.txt", Speedmem);
	 $readmemh("CoverArt/Pause.txt", Pausemem);
	 $readmemh("CoverArt/Play.txt", Playmem);
	 $readmemh("CoverArt/GrenadeTitle.txt", Titlemem);
	 $readmemh("CoverArt/JustTitle.txt", Title2mem);
end

always_ff @ (posedge CLOCK) begin
	if (SecondSong) 
		CoverArtColor<= JustArtmem[CoverPixel];
	else
		CoverArtColor<= GrenadeArtmem[CoverPixel];

	if (RW)
		PlayPauseColor<= Playmem[PlayPausePixel];
	else
		PlayPauseColor<= Pausemem[PlayPausePixel];

	if (SecondSong) 
		TitleColor<= Title2mem[TitlePixel];
	else
		TitleColor<= Titlemem[TitlePixel];

	SpeedColor<= Speedmem[SpeedPixel];
	
end
endmodule
